module vulkan

#flag -I $env('VULKAN_SDK')/Include
#flag -L $env('VULKAN_SDK')/Libs
#flag -lvulkan-1