module vulkan

#flag -lvulkan